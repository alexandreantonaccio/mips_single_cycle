`timescale 1ns/1ps

module bne_cpu_tb();

    logic clk, reset;
    logic [31:0] writedata, dataadr;
    logic memwrite;
    
    // Instanciação da CPU
    bne_cpu dut (
        .clk(clk),
        .reset(reset),
        .writedata(writedata),
        .dataadr(dataadr),
        .memwrite(memwrite)
    );
    
    // Gerador de clock (período 10ns)
    always begin
        clk = 1; #5;
        clk = 0; #5;
    end
    
    // Inicialização e sequência de teste
    initial begin
        // Inicializa registros e memórias
        reset = 1;
        #10; 
        reset = 0;
        
        // Aguarda execução completa (ajustar conforme necessidade)
        #1000;
        
        $finish;
    end
    initial begin
		  forever @(negedge clk) begin
			 if (!reset) begin
				$display("t0=%h t1=%h t2=%h t3=%h t4=%h t5=%h t6=%h t7=%h",
							dut.cpu.dp.rf.rf[8],  // $t0
							dut.cpu.dp.rf.rf[9],  // $t1
							dut.cpu.dp.rf.rf[10], // $t2
							dut.cpu.dp.rf.rf[11], // $t3
							dut.cpu.dp.rf.rf[12], // $t4
							dut.cpu.dp.rf.rf[13], // $t5
							dut.cpu.dp.rf.rf[14], // $t6
							dut.cpu.dp.rf.rf[15]);// $t7
							
			 end
		  end
		end

    initial begin
        $display("Tempo\t PC       \t Instr\t\t Operação\t Reg/Mem\t Dados");
        $display("------------------------------------------------------------------");
        
        // Formatação personalizada para visualização
        forever @(negedge clk) begin
            if (!reset) begin
                $write("%4d:\t %h\t %h\t", $time, dut.pc, dut.instr);
                
                // Decodificação básica para exibição
                casez (dut.instr[31:26])
                    6'b000000: $write("R-type\t\t");
                    6'b100011: $write("LW    \t\t");
                    6'b101011: $write("SW    \t\t");
                    6'b000100: $write("BEQ   \t\t");
                    6'b000101: $write("BNE   \t\t");
                    6'b001000: $write("ADDI  \t\t");
                    6'b000010: $write("J     \t\t");
                    default:   $write("Unknown\t\t");
                endcase
                
                if (memwrite) begin
                    $write("Mem[%h] = %h", dataadr, writedata);
                end
                $display();
            end
        end
    end
endmodule